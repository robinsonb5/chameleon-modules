library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------

entity chameleon_mergeinputs is
	generic (
		joybits : integer :=8;
		button1 : integer :=4;
		button2 : integer :=5;
		button3 : integer :=6;
		button4 : integer :=7
	);
	port (
		clk : in std_logic; -- 100 MHz input clock
		reset_n : in std_logic;
		ena_1mhz : in std_logic;
		ir_data : in std_logic;
		button_menu_n : in std_logic;
		c64_joy1 : in unsigned(6 downto 0);
		c64_joy2 : in unsigned(6 downto 0);
		c64_joy3 : in unsigned(6 downto 0);
		c64_joy4 : in unsigned(6 downto 0);
		c64_keys : in unsigned(63 downto 0);
		c64_joykey_ena : in std_logic;

		joy1_out : out unsigned(joybits-1 downto 0);
		joy2_out : out unsigned(joybits-1 downto 0);
		joy3_out : out unsigned(joybits-1 downto 0);
		joy4_out : out unsigned(joybits-1 downto 0);
		menu_out_n : out std_logic
	);
end entity;

architecture rtl of chameleon_mergeinputs is

-- CDTV pad signals:
signal ir : std_logic;
signal ir_d : std_logic;
signal cdtv_port : std_logic;
signal cdtv_joya : unsigned(5 downto 0);
signal cdtv_joyb : unsigned(5 downto 0);
signal cdtv_power : std_logic;
signal cdtv_play : std_logic;
signal cdtv_volup : std_logic;
signal cdtv_voldown : std_logic;

-- c64 keyboard-related signals
signal keys_safe : std_logic;
signal c64_menu : std_logic :='1';
signal c64_start1 : std_logic :='1';
signal c64_select1 :std_logic :='1';
signal c64_start2 : std_logic :='1';
signal c64_select2 : std_logic :='1';

-- Merged signals for buttons 3/4	
signal porta_start : std_logic;
signal porta_select : std_logic;
signal portb_start : std_logic;
signal portb_select : std_logic;

begin

	-- Synchronise IR signal
	process (clk)
	begin
		if rising_edge(clk) then
			ir_d<=ir_data;
			ir<=ir_d;
		end if;
	end process;


	cdtv : entity work.chameleon_cdtv_remote
	port map(
		clk => clk,
		ena_1mhz => ena_1mhz,
		ir => ir,
		key_power => cdtv_power,
		key_play => cdtv_play,
		joystick_a => cdtv_joya,
		joystick_b => cdtv_joyb,
		key_vol_up => cdtv_volup,
		key_vol_dn => cdtv_voldown,
		currentport => cdtv_port
	);

	keys_safe <= '1' when c64_joy1="1111111" else '0';

	-- Update c64 keys only when the joystick isn't active.
	process (clk,reset_n)
	begin
		if reset_n='0' then
			c64_start1<='1';
			c64_select1<='1';
			c64_start2<='1';
			c64_select2<='1';
			c64_menu<='1';
		elsif rising_edge(clk) then
			if keys_safe='1' then
				c64_start1 <= not c64_joykey_ena or c64_keys(8); -- Return
				c64_select1 <= not c64_joykey_ena or c64_keys(38); -- Right shift
				c64_start2 <= not c64_joykey_ena or c64_keys(63); -- Run/stop
				c64_select2 <= not c64_joykey_ena or c64_keys(57); -- Left shift;
				c64_menu <= not c64_joykey_ena or c64_keys(15); -- Left arrow;
			end if;
		end if;
	end process;

	-- 3rd and 4th buttons, active low
	porta_start <= (cdtv_port or not cdtv_play) and c64_start1;
	porta_select <= ((cdtv_port or not cdtv_volup) and c64_select1) and c64_joy1(6);

	portb_start <= (not cdtv_port or not cdtv_play) and c64_start2;
	portb_select <= ((not cdtv_port or not cdtv_volup) and c64_select2) and c64_joy2(6);

	-- Output mapping
	process(c64_joy1,c64_joy2,c64_joy3,c64_joy4,cdtv_joya,cdtv_joyb,porta_select,portb_select,porta_start,portb_start)
	begin
		joy1_out<=(others=>'1');
		joy2_out<=(others=>'1');
		joy3_out<=(others=>'1');
		joy4_out<=(others=>'1');

		joy1_out(3 downto 0)<=c64_joy1(3 downto 0) and cdtv_joya(3 downto 0);
		joy2_out(3 downto 0)<=c64_joy2(3 downto 0) and cdtv_joyb(3 downto 0);
		joy3_out(3 downto 0)<=c64_joy3(3 downto 0);
		joy4_out(3 downto 0)<=c64_joy4(3 downto 0);

		-- First button
		joy1_out(button1)<=c64_joy1(4) and cdtv_joya(4);
		joy2_out(button1)<=c64_joy2(4) and cdtv_joyb(4);
		joy3_out(button1)<=c64_joy3(4);
		joy4_out(button1)<=c64_joy4(4);

		-- Second button
		joy1_out(button2)<=c64_joy1(5) and cdtv_joya(5);
		joy2_out(button2)<=c64_joy2(5) and cdtv_joyb(5);
		joy3_out(button2)<=c64_joy3(5);
		joy4_out(button2)<=c64_joy4(5);

		-- Third button
		joy1_out(button3)<=porta_select and c64_joy1(6);
		joy2_out(button3)<=portb_select and c64_joy2(6);
		joy3_out(button3)<=c64_joy3(6);
		joy4_out(button3)<=c64_joy4(6);

		-- Fourth button
		joy1_out(button4)<=porta_start;
		joy2_out(button4)<=portb_start;
		joy3_out(button4)<='1';
		joy4_out(button4)<='1';
	end process;

	menu_out_n<=button_menu_n and c64_menu and not cdtv_power;
	
end architecture;
